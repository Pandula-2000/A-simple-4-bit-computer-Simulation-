CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 70 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
68
13 Logic Switch~
5 568 759 0 1 11
0 12
0
0 0 20576 0
2 0V
-6 -16 8 -8
3 V28
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6118 0 0
2
44470.6 17
0
13 Logic Switch~
5 590 768 0 1 11
0 13
0
0 0 20576 0
2 0V
-6 -16 8 -8
3 V29
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
34 0 0
2
44470.6 16
0
13 Logic Switch~
5 691 804 0 1 11
0 17
0
0 0 20576 0
2 0V
-6 -16 8 -8
3 V30
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6357 0 0
2
44470.6 15
0
13 Logic Switch~
5 667 795 0 1 11
0 14
0
0 0 20576 0
2 0V
-6 -16 8 -8
3 V31
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
319 0 0
2
44470.6 14
0
13 Logic Switch~
5 612 777 0 1 11
0 16
0
0 0 20576 0
2 0V
-6 -16 8 -8
3 V32
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3976 0 0
2
44470.6 13
0
13 Logic Switch~
5 638 786 0 1 11
0 15
0
0 0 20576 0
2 0V
-6 -16 8 -8
3 V33
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7634 0 0
2
44470.6 12
0
13 Logic Switch~
5 784 840 0 1 11
0 21
0
0 0 20576 0
2 0V
-6 -16 8 -8
3 V34
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
523 0 0
2
44470.6 11
0
13 Logic Switch~
5 761 831 0 1 11
0 18
0
0 0 20576 0
2 0V
-6 -16 8 -8
3 V35
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6748 0 0
2
44470.6 10
0
13 Logic Switch~
5 713 813 0 1 11
0 20
0
0 0 20576 0
2 0V
-6 -16 8 -8
3 V36
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6901 0 0
2
44470.6 9
0
13 Logic Switch~
5 737 822 0 1 11
0 19
0
0 0 20576 0
2 0V
-6 -16 8 -8
3 V37
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
842 0 0
2
44470.6 8
0
13 Logic Switch~
5 844 941 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 20704 0
2 5V
-6 -16 8 -8
3 V38
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3277 0 0
2
44470.6 7
0
13 Logic Switch~
5 847 897 0 1 11
0 24
0
0 0 20576 0
2 0V
-6 -16 8 -8
3 V39
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4212 0 0
2
44470.6 6
0
13 Logic Switch~
5 1020 611 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 20704 0
2 5V
-6 -16 8 -8
3 V45
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4720 0 0
2
44470.6 5
0
13 Logic Switch~
5 1150 951 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 20576 180
2 5V
-6 -16 8 -8
3 V46
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5551 0 0
2
44470.6 0
0
13 Logic Switch~
5 1007 541 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 20720 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6986 0 0
2
44470.5 0
0
13 Logic Switch~
5 646 447 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 20720 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8745 0 0
2
44470.5 0
0
13 Logic Switch~
5 445 527 0 1 11
0 68
0
0 0 20720 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9592 0 0
2
44470.5 0
0
13 Logic Switch~
5 454 814 0 1 11
0 73
0
0 0 20720 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8748 0 0
2
44470.5 1
0
13 Logic Switch~
5 453 784 0 1 11
0 74
0
0 0 20720 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7168 0 0
2
44470.5 2
0
13 Logic Switch~
5 444 683 0 1 11
0 42
0
0 0 20720 0
2 0V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
631 0 0
2
44470.5 3
0
13 Logic Switch~
5 449 749 0 1 11
0 75
0
0 0 20720 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9466 0 0
2
44470.5 4
0
13 Logic Switch~
5 449 625 0 1 11
0 72
0
0 0 20720 0
2 0V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3266 0 0
2
44470.5 5
0
13 Logic Switch~
5 447 604 0 1 11
0 71
0
0 0 20720 0
2 0V
-6 -16 8 -8
3 V14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7693 0 0
2
44470.5 6
0
13 Logic Switch~
5 445 581 0 1 11
0 66
0
0 0 20720 0
2 0V
-6 -16 8 -8
3 V15
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3723 0 0
2
44470.5 7
0
13 Logic Switch~
5 444 558 0 1 11
0 67
0
0 0 20720 0
2 0V
-6 -16 8 -8
3 V16
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3440 0 0
2
44470.5 8
0
13 Logic Switch~
5 472 209 0 1 11
0 62
0
0 0 20592 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6263 0 0
2
5.90002e-315 0
0
13 Logic Switch~
5 446 200 0 1 11
0 63
0
0 0 20592 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4900 0 0
2
5.90002e-315 5.26354e-315
0
13 Logic Switch~
5 392 182 0 1 11
0 65
0
0 0 20592 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8783 0 0
2
5.90002e-315 5.30499e-315
0
13 Logic Switch~
5 419 191 0 1 11
0 64
0
0 0 20592 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3221 0 0
2
5.90002e-315 5.32571e-315
0
7 74LS244
143 1084 740 0 18 37
0 8 9 10 7 76 77 78 79 6
5 4 3 80 81 82 83 22 84
0
0 0 4832 0
7 74LS244
-24 -60 25 -52
3 U15
-10 -61 11 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP14
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 512 1 0 0 0
1 U
3215 0 0
2
44470.6 24
0
6 1K RAM
79 870 795 0 20 41
0 12 13 16 15 14 17 20 19 18
21 85 86 87 88 8 9 10 7 24
11
0
0 0 4832 0
5 RAM1K
-17 -19 18 -11
3 U16
-11 -70 10 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
7903 0 0
2
44470.6 23
0
7 74LS244
143 1087 866 0 18 37
0 6 5 4 3 89 90 91 92 8
9 10 7 93 94 95 96 23 97
0
0 0 4832 180
7 74LS244
-24 -60 25 -52
3 U17
-17 -61 4 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP14
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 512 1 0 0 0
1 U
7121 0 0
2
44470.6 18
0
7 74LS244
143 1107 172 0 18 37
0 98 99 100 101 41 40 39 38 102
103 104 105 3 4 5 6 106 25
0
0 0 4848 180
7 74LS244
-24 -60 25 -52
2 U6
-13 -61 1 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP14
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 512 1 0 0 0
1 U
4484 0 0
2
44470.5 0
0
7 74LS273
150 1034 457 0 18 37
0 35 34 107 108 109 110 6 5 4
3 111 112 113 114 26 27 28 29
0
0 0 4848 180
7 74LS273
-24 -60 25 -52
2 U3
-13 -61 1 -53
0
16 DVCC=20;DGND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
5996 0 0
2
5.90002e-315 0
0
7 74LS273
150 728 384 0 18 37
0 37 36 115 116 117 118 6 5 4
3 119 120 121 122 30 31 32 33
0
0 0 4848 0
7 74LS273
-24 -60 25 -52
2 U8
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
7804 0 0
2
5.90002e-315 0
0
9 Inverter~
13 1660 649 0 2 22
0 41 48
0
0 0 112 180
6 74LS04
-21 -19 21 -11
3 U7F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
5523 0 0
2
5.90002e-315 5.34643e-315
0
9 Inverter~
13 1618 406 0 2 22
0 46 43
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U7B
20 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3330 0 0
2
5.90002e-315 5.3568e-315
0
9 2-In AND~
219 1541 614 0 3 22
0 44 43 45
0
0 0 112 180
6 74LS08
-21 -24 21 -16
3 U9C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3465 0 0
2
5.90002e-315 5.36716e-315
0
9 2-In AND~
219 1541 537 0 3 22
0 38 42 47
0
0 0 112 180
6 74LS08
-21 -24 21 -16
3 U9D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
8396 0 0
2
5.90002e-315 5.37752e-315
0
14 Logic Display~
6 1469 544 0 1 2
10 46
0
0 0 53360 90
6 100MEG
3 -16 45 -8
2 L5
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3685 0 0
2
5.90002e-315 5.38788e-315
0
14 Logic Display~
6 1471 577 0 1 2
10 47
0
0 0 53360 90
6 100MEG
3 -16 45 -8
2 L6
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7849 0 0
2
5.90002e-315 5.39306e-315
0
14 Logic Display~
6 1474 608 0 1 2
10 45
0
0 0 53360 90
6 100MEG
3 -16 45 -8
2 L7
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6343 0 0
2
5.90002e-315 5.39824e-315
0
9 Inverter~
13 1656 564 0 2 22
0 38 51
0
0 0 112 180
6 74LS04
-21 -19 21 -11
3 U7C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
7376 0 0
2
5.90002e-315 5.40342e-315
0
9 Inverter~
13 1656 591 0 2 22
0 39 50
0
0 0 112 180
6 74LS04
-21 -19 21 -11
3 U7D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
9156 0 0
2
5.90002e-315 5.4086e-315
0
9 Inverter~
13 1660 616 0 2 22
0 40 49
0
0 0 112 180
6 74LS04
-21 -19 21 -11
3 U7E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
5776 0 0
2
5.90002e-315 5.41378e-315
0
9 4-In AND~
219 1607 614 0 5 22
0 48 49 50 51 44
0
0 0 624 180
6 74LS21
-21 -28 21 -20
4 U10A
-16 -28 12 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 4 0
1 U
7207 0 0
2
5.90002e-315 5.41896e-315
0
14 Logic Display~
6 1545 237 0 1 2
10 38
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4459 0 0
2
5.90002e-315 5.42414e-315
0
14 Logic Display~
6 1575 234 0 1 2
10 39
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3760 0 0
2
5.90002e-315 5.42933e-315
0
14 Logic Display~
6 1607 235 0 1 2
10 40
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
754 0 0
2
5.90002e-315 5.43192e-315
0
14 Logic Display~
6 1633 235 0 1 2
10 41
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9767 0 0
2
5.90002e-315 5.43451e-315
0
6 74136~
219 1287 352 0 3 22
0 26 42 55
0
0 0 112 0
7 74LS136
-24 -24 25 -16
4 U11A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7978 0 0
2
5.90002e-315 5.4371e-315
0
6 74136~
219 1283 393 0 3 22
0 27 42 54
0
0 0 112 0
7 74LS136
-24 -24 25 -16
4 U11B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3142 0 0
2
5.90002e-315 5.43969e-315
0
6 74136~
219 1287 431 0 3 22
0 28 42 53
0
0 0 112 0
7 74LS136
-24 -24 25 -16
4 U11C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3284 0 0
2
5.90002e-315 5.44228e-315
0
6 74136~
219 1284 470 0 3 22
0 29 42 52
0
0 0 112 0
7 74LS136
-24 -24 25 -16
4 U11D
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
659 0 0
2
5.90002e-315 5.44487e-315
0
7 74LS283
152 1497 303 0 14 29
0 30 31 32 33 55 54 53 52 42
38 39 40 41 46
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
3 U13
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 0 1 0 0 0
1 U
3800 0 0
2
5.90002e-315 5.44746e-315
0
9 2-In AND~
219 940 506 0 3 22
0 66 68 34
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6792 0 0
2
44470.5 9
0
9 2-In AND~
219 604 498 0 3 22
0 67 68 36
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3701 0 0
2
44470.5 10
0
9 Inverter~
13 597 603 0 2 22
0 71 70
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
6316 0 0
2
44470.5 13
0
9 Inverter~
13 511 625 0 2 22
0 72 69
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U5F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
8734 0 0
2
44470.5 14
0
9 Inverter~
13 478 813 0 2 22
0 73 25
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U5E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
7988 0 0
2
44470.5 15
0
9 Inverter~
13 478 783 0 2 22
0 74 60
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U5D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3217 0 0
2
44470.5 16
0
9 Inverter~
13 473 749 0 2 22
0 75 61
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U5C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3965 0 0
2
44470.5 17
0
7 74LS244
143 873 368 0 18 37
0 30 31 32 33 26 27 28 29 6
5 4 3 6 5 4 3 70 69
0
0 0 4848 90
7 74LS244
-24 -60 25 -52
2 U4
54 -6 68 2
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP14
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 0 1 0 0 0
1 U
8239 0 0
2
44470.5 18
0
14 Logic Display~
6 908 53 0 1 2
10 56
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
828 0 0
2
5.90002e-315 5.45005e-315
0
14 Logic Display~
6 884 54 0 1 2
10 57
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6187 0 0
2
5.90002e-315 5.45264e-315
0
14 Logic Display~
6 860 56 0 1 2
10 58
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7107 0 0
2
5.90002e-315 5.45523e-315
0
14 Logic Display~
6 836 57 0 1 2
10 59
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6433 0 0
2
5.90002e-315 5.45782e-315
0
7 74LS244
143 718 164 0 18 37
0 6 5 4 3 65 64 63 62 59
58 57 56 6 5 4 3 60 61
0
0 0 4848 0
7 74LS244
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP14
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 0 1 0 0 0
1 U
8559 0 0
2
5.90002e-315 5.463e-315
0
157
4 0 3 0 0 4096 0 32 0 0 8 2
1113 870
1191 870
3 0 4 0 0 4096 0 32 0 0 9 2
1113 879
1181 879
2 0 5 0 0 4096 0 32 0 0 10 2
1113 888
1173 888
9 0 6 0 0 4096 0 30 0 0 11 2
1116 713
1163 713
10 0 5 0 0 0 0 30 0 0 10 2
1116 722
1173 722
11 0 4 0 0 0 0 30 0 0 9 2
1116 731
1181 731
12 0 3 0 0 0 0 30 0 0 8 2
1116 740
1191 740
0 0 3 0 0 4096 0 0 0 70 0 2
1191 295
1191 892
0 0 4 0 0 4096 0 0 0 71 0 2
1181 285
1181 893
0 0 5 0 0 4096 0 0 0 72 0 2
1173 273
1173 896
0 1 6 0 0 4096 0 0 32 73 0 3
1163 264
1163 897
1113 897
18 0 7 0 0 4096 0 31 0 0 38 2
902 840
977 840
0 15 8 0 0 4096 0 0 31 37 0 2
953 813
902 813
0 16 9 0 0 4096 0 0 31 40 0 2
962 822
902 822
0 17 10 0 0 4096 0 0 31 39 0 2
969 831
902 831
20 1 11 0 0 8320 0 31 11 0 0 4
908 768
912 768
912 941
856 941
1 1 12 0 0 8320 0 1 31 0 0 2
580 759
838 759
2 1 13 0 0 4224 0 31 2 0 0 2
838 768
602 768
5 1 14 0 0 4224 0 31 4 0 0 2
838 795
679 795
4 1 15 0 0 4240 0 31 6 0 0 2
838 786
650 786
3 1 16 0 0 4224 0 31 5 0 0 2
838 777
624 777
1 6 17 0 0 4224 0 3 31 0 0 2
703 804
838 804
9 1 18 0 0 12416 0 31 8 0 0 2
838 831
773 831
8 1 19 0 0 4224 0 31 10 0 0 2
838 822
749 822
7 1 20 0 0 4224 0 31 9 0 0 2
838 813
725 813
1 10 21 0 0 12416 0 7 31 0 0 2
796 840
838 840
17 1 22 0 0 8320 0 30 13 0 0 3
1046 704
1032 704
1032 611
17 1 23 0 0 8320 0 32 14 0 0 4
1119 906
1134 906
1134 951
1136 951
9 0 8 0 0 4096 0 32 0 0 37 2
1049 897
953 897
10 0 9 0 0 4096 0 32 0 0 40 2
1049 888
962 888
11 0 10 0 0 4096 0 32 0 0 39 2
1049 879
969 879
12 0 7 0 0 0 0 32 0 0 38 2
1049 870
977 870
1 0 8 0 0 4096 0 30 0 0 37 2
1052 713
953 713
2 0 9 0 0 4096 0 30 0 0 40 2
1052 722
962 722
3 0 10 0 0 4096 0 30 0 0 39 2
1052 731
969 731
4 0 7 0 0 0 0 30 0 0 38 2
1052 740
977 740
0 0 8 0 0 4224 0 0 0 0 0 2
953 680
953 919
0 0 7 0 0 4224 0 0 0 0 0 2
977 681
977 918
0 0 10 0 0 4224 0 0 0 0 0 2
969 680
969 920
0 0 9 0 0 4224 0 0 0 0 0 2
962 679
962 921
1 0 24 0 0 4096 0 12 0 0 42 2
859 897
859 896
19 1 24 0 0 8320 0 31 0 0 0 6
908 759
916 759
916 907
864 907
864 896
855 896
18 0 25 0 0 4096 0 33 0 0 76 3
1139 167
1211 167
1211 176
0 5 26 0 0 4096 0 0 63 63 0 3
949 442
886 442
886 399
0 6 27 0 0 4096 0 0 63 62 0 3
956 434
895 434
895 399
0 7 28 0 0 4096 0 0 63 61 0 3
964 423
904 423
904 399
0 8 29 0 0 4096 0 0 63 60 0 3
970 416
913 416
913 399
7 0 6 0 0 0 0 34 0 0 73 3
1060 443
1104 443
1104 264
8 0 5 0 0 0 0 34 0 0 72 3
1060 434
1116 434
1116 273
9 0 4 0 0 0 0 34 0 0 71 3
1060 425
1128 425
1128 285
10 0 3 0 0 0 0 34 0 0 70 3
1060 416
1137 416
1137 295
0 1 30 0 0 4096 0 0 63 67 0 3
780 402
841 402
841 399
0 2 31 0 0 4096 0 0 63 66 0 3
788 411
850 411
850 399
0 3 32 0 0 4096 0 0 63 65 0 3
798 420
859 420
859 399
18 4 33 0 0 8320 0 35 63 0 0 4
760 429
760 436
868 436
868 399
9 0 4 0 0 0 0 35 0 0 71 3
696 420
628 420
628 285
7 0 6 0 0 0 0 35 0 0 73 3
696 402
606 402
606 264
8 0 5 0 0 0 0 35 0 0 72 3
696 411
617 411
617 273
10 0 3 0 0 0 0 35 0 0 70 3
696 429
641 429
641 295
1 18 29 0 0 12416 0 54 34 0 0 6
1268 461
1180 461
1180 369
970 369
970 416
996 416
1 17 28 0 0 12416 0 53 34 0 0 7
1271 422
1191 422
1191 357
964 357
964 424
996 424
996 425
1 16 27 0 0 12416 0 52 34 0 0 6
1267 384
1209 384
1209 350
956 350
956 434
996 434
1 15 26 0 0 4224 0 51 34 0 0 5
1271 343
949 343
949 442
996 442
996 443
0 4 33 0 0 8320 0 0 55 55 0 5
810 436
810 327
1273 327
1273 294
1465 294
17 3 32 0 0 12416 0 35 55 0 0 6
760 420
798 420
798 323
1268 323
1268 285
1465 285
16 2 31 0 0 12416 0 35 55 0 0 6
760 411
788 411
788 318
1263 318
1263 276
1465 276
15 1 30 0 0 12416 0 35 55 0 0 6
760 402
780 402
780 313
1256 313
1256 267
1465 267
3 2 34 0 0 12416 0 56 34 0 0 6
961 506
983 506
983 515
1117 515
1117 488
1060 488
1 1 35 0 0 8320 0 34 15 0 0 4
1066 497
1066 543
1019 543
1019 541
0 0 3 0 0 4224 0 0 0 0 0 2
590 295
1224 295
0 0 4 0 0 4224 0 0 0 0 0 2
590 285
1224 285
0 0 5 0 0 4224 0 0 0 0 0 2
588 273
1227 273
0 0 6 0 0 4224 0 0 0 0 0 2
590 264
1229 264
2 3 36 0 0 8320 0 35 57 0 0 4
696 357
680 357
680 498
625 498
1 1 37 0 0 8320 0 16 35 0 0 4
658 447
659 447
659 348
690 348
2 0 25 0 0 12416 0 60 0 0 43 7
499 813
512 813
512 667
1084 667
1084 238
1211 238
1211 172
16 0 6 0 0 0 0 33 0 0 73 4
1069 131
1069 130
991 130
991 264
15 0 5 0 0 0 0 33 0 0 72 4
1069 140
1069 139
1005 139
1005 273
14 0 4 0 0 0 0 33 0 0 71 4
1069 149
1069 148
1023 148
1023 285
13 0 3 0 0 0 0 33 0 0 70 4
1069 158
1069 157
1034 157
1034 295
0 8 38 0 0 8320 0 0 33 112 0 4
1756 294
1756 130
1133 130
1133 131
7 0 39 0 0 8320 0 33 0 0 111 4
1133 140
1133 139
1766 139
1766 303
0 6 40 0 0 8320 0 0 33 110 0 4
1776 312
1776 148
1133 148
1133 149
5 0 41 0 0 8320 0 33 0 0 109 4
1133 158
1133 157
1784 157
1784 321
2 0 42 0 0 4096 0 53 0 0 87 2
1271 440
1222 440
2 0 42 0 0 0 0 52 0 0 87 2
1267 402
1222 402
1 2 42 0 0 16512 0 20 51 0 0 7
456 683
456 646
643 646
643 644
1222 644
1222 361
1271 361
2 0 43 0 0 8192 0 37 0 0 89 3
1621 424
1620 424
1620 445
2 0 43 0 0 24704 0 38 0 0 0 7
1559 605
1571 605
1571 570
1613 570
1613 517
1620 517
1620 440
1 5 44 0 0 4224 0 38 46 0 0 3
1559 623
1580 623
1580 614
1 3 45 0 0 8320 0 42 38 0 0 3
1489 611
1489 614
1514 614
0 1 46 0 0 4096 0 0 37 97 0 3
1529 369
1621 369
1621 388
1 0 41 0 0 0 0 50 0 0 109 2
1633 253
1633 321
1 0 40 0 0 0 0 49 0 0 110 2
1607 253
1607 312
1 0 39 0 0 0 0 48 0 0 111 2
1575 252
1575 303
1 0 38 0 0 0 0 47 0 0 112 2
1545 255
1545 294
1 14 46 0 0 8320 0 40 55 0 0 5
1484 547
1506 547
1506 405
1529 405
1529 348
1 3 47 0 0 8320 0 41 39 0 0 3
1486 580
1514 580
1514 537
0 1 38 0 0 0 0 0 39 112 0 3
1585 294
1585 546
1559 546
0 2 42 0 0 0 0 0 39 113 0 4
1454 451
1577 451
1577 528
1559 528
0 1 41 0 0 0 0 0 36 109 0 4
1715 321
1715 650
1681 650
1681 649
1 0 40 0 0 0 0 45 0 0 110 3
1681 616
1702 616
1702 312
0 1 39 0 0 0 0 0 44 111 0 3
1687 303
1687 591
1677 591
1 0 38 0 0 0 0 43 0 0 112 3
1677 564
1675 564
1675 294
1 2 48 0 0 4224 0 46 36 0 0 4
1625 627
1625 650
1645 650
1645 649
2 2 49 0 0 8320 0 45 46 0 0 3
1645 616
1645 618
1625 618
2 3 50 0 0 8320 0 44 46 0 0 4
1641 591
1634 591
1634 609
1625 609
2 4 51 0 0 8320 0 43 46 0 0 3
1641 564
1625 564
1625 600
13 0 41 0 0 0 0 55 0 0 0 2
1529 321
1795 321
12 0 40 0 0 0 0 55 0 0 0 2
1529 312
1800 312
11 0 39 0 0 0 0 55 0 0 0 2
1529 303
1790 303
10 0 38 0 0 0 0 55 0 0 0 2
1529 294
1796 294
0 9 42 0 0 0 0 0 55 87 0 4
1222 492
1454 492
1454 348
1465 348
2 0 42 0 0 0 0 54 0 0 87 2
1268 479
1222 479
3 8 52 0 0 8320 0 54 55 0 0 5
1317 470
1438 470
1438 329
1465 329
1465 330
3 7 53 0 0 8320 0 53 55 0 0 5
1320 431
1425 431
1425 320
1465 320
1465 321
3 6 54 0 0 4224 0 52 55 0 0 5
1316 393
1412 393
1412 311
1465 311
1465 312
3 5 55 0 0 4224 0 51 55 0 0 5
1320 352
1400 352
1400 302
1465 302
1465 303
13 0 6 0 0 0 0 68 0 0 73 3
750 182
758 182
758 264
14 0 5 0 0 0 0 68 0 0 72 3
750 191
765 191
765 273
15 0 4 0 0 0 0 68 0 0 71 3
750 200
773 200
773 285
16 0 3 0 0 0 0 68 0 0 70 3
750 209
780 209
780 295
12 1 56 0 0 4224 0 68 64 0 0 3
750 164
908 164
908 71
11 1 57 0 0 4224 0 68 65 0 0 3
750 155
884 155
884 72
10 1 58 0 0 4224 0 68 66 0 0 3
750 146
860 146
860 74
9 1 59 0 0 4224 0 68 67 0 0 3
750 137
836 137
836 75
17 2 60 0 0 8320 0 68 61 0 0 6
680 128
548 128
548 660
503 660
503 783
499 783
1 0 6 0 0 0 0 68 0 0 73 3
686 137
648 137
648 264
2 0 5 0 0 0 0 68 0 0 72 3
686 146
657 146
657 273
3 0 4 0 0 0 0 68 0 0 71 3
686 155
667 155
667 285
4 0 3 0 0 0 0 68 0 0 70 3
686 164
677 164
677 295
2 18 61 0 0 12416 0 62 68 0 0 5
494 749
494 652
517 652
517 173
680 173
1 0 62 0 0 4096 0 26 0 0 134 2
484 209
502 209
8 0 62 0 0 4224 0 68 0 0 0 2
686 209
499 209
7 1 63 0 0 4224 0 68 27 0 0 2
686 200
458 200
6 1 64 0 0 4224 0 68 29 0 0 2
686 191
431 191
5 1 65 0 0 4224 0 68 28 0 0 2
686 182
404 182
1 1 66 0 0 4224 0 24 56 0 0 4
457 581
893 581
893 497
916 497
1 1 67 0 0 4224 0 25 57 0 0 4
456 558
555 558
555 489
580 489
2 0 68 0 0 8192 0 56 0 0 142 3
916 515
905 515
905 527
2 0 68 0 0 8192 0 57 0 0 142 3
580 507
566 507
566 527
1 0 68 0 0 4224 0 17 0 0 0 2
457 527
917 527
18 2 69 0 0 8320 0 63 59 0 0 3
877 405
877 625
532 625
17 2 70 0 0 8320 0 63 58 0 0 3
832 405
832 603
618 603
1 1 71 0 0 4224 0 58 23 0 0 4
582 603
474 603
474 604
459 604
1 1 72 0 0 4224 0 59 22 0 0 2
496 625
461 625
1 1 73 0 0 8320 0 60 18 0 0 3
463 813
463 814
466 814
1 1 74 0 0 8320 0 61 19 0 0 3
463 783
463 784
465 784
1 1 75 0 0 4224 0 62 21 0 0 2
458 749
461 749
13 0 6 0 0 0 0 63 0 0 73 2
886 335
886 264
14 0 5 0 0 0 0 63 0 0 72 2
895 335
895 273
15 0 4 0 0 0 0 63 0 0 71 2
904 335
904 285
16 0 3 0 0 0 0 63 0 0 70 2
913 335
913 295
9 0 6 0 0 0 0 63 0 0 73 2
841 335
841 264
10 0 5 0 0 0 0 63 0 0 72 2
850 335
850 273
11 0 4 0 0 0 0 63 0 0 71 2
859 335
859 285
12 0 3 0 0 0 0 63 0 0 70 2
868 335
868 295
23
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
746 881 845 896
760 892 830 903
10 RAM ENABLE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
357 176 392 200
368 185 380 201
2 x3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
380 186 415 210
391 195 403 211
2 x2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
407 196 442 220
418 204 430 220
2 x1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
437 208 472 232
448 217 460 233
2 x0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
630 717 695 741
641 726 683 742
7 ADDRESS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
1156 924 1221 968
1167 933 1209 965
18 RAM=BUS 
(WRITE)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
951 582 1016 626
962 591 1004 623
16 RAM=BUS
(READ)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
747 925 830 949
758 934 818 950
10 READ/WRITE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
392 513 433 534
400 520 424 535
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
326 800 441 821
335 807 431 822
12 DBUS=ALU_OUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
373 769 438 790
381 776 429 791
6 Z=DBUS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
369 734 434 755
377 741 425 756
6 DBUS=X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
362 676 427 700
373 685 415 701
7 SUB '1'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
367 656 426 680
375 665 417 681
7 ADD '0'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
358 615 425 636
367 621 415 636
6 DBUS=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
359 591 426 612
368 597 416 612
6 DBUS=A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
354 568 427 589
362 574 418 589
7 B<<DBUS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
355 546 428 567
363 553 419 568
7 A<<DBUS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1673 263 1749 286
1686 273 1735 288
7 ALU_OUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1422 532 1457 553
1431 539 1447 554
2 CF
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1423 597 1458 618
1432 603 1448 618
2 ZF
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1422 564 1457 585
1431 571 1447 586
2 NF
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
